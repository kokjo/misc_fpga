module font_8x8 (clk, rst, ch, bitmap);
    input clk; input rst;
    input [7:0] ch;
    output reg [63:0] bitmap;
    reg [63:0] font [0:127];

    initial begin
        font[8'h00] = 64'h0000000000000000;
        font[8'h01] = 64'h0000000000000000;
        font[8'h02] = 64'h0000000000000000;
        font[8'h03] = 64'h0000000000000000;
        font[8'h04] = 64'h0000000000000000;
        font[8'h05] = 64'h0000000000000000;
        font[8'h06] = 64'h0000000000000000;
        font[8'h07] = 64'h0000000000000000;
        font[8'h08] = 64'h0000000000000000;
        font[8'h09] = 64'h0000000000000000;
        font[8'h0a] = 64'h0000000000000000;
        font[8'h0b] = 64'h0000000000000000;
        font[8'h0c] = 64'h0000000000000000;
        font[8'h0d] = 64'h0000000000000000;
        font[8'h0e] = 64'h0000000000000000;
        font[8'h0f] = 64'h0000000000000000;
        font[8'h10] = 64'h0000000000000000;
        font[8'h11] = 64'h0000000000000000;
        font[8'h12] = 64'h0000000000000000;
        font[8'h13] = 64'h0000000000000000;
        font[8'h14] = 64'h0000000000000000;
        font[8'h15] = 64'h0000000000000000;
        font[8'h16] = 64'h0000000000000000;
        font[8'h17] = 64'h0000000000000000;
        font[8'h18] = 64'h0000000000000000;
        font[8'h19] = 64'h0000000000000000;
        font[8'h1a] = 64'h0000000000000000;
        font[8'h1b] = 64'h0000000000000000;
        font[8'h1c] = 64'h0000000000000000;
        font[8'h1d] = 64'h0000000000000000;
        font[8'h1e] = 64'h0000000000000000;
        font[8'h1f] = 64'h0000000000000000;
        font[8'h20] = 64'h0000000000000000;
        font[8'h21] = 64'h183C3C1818001800;
        font[8'h22] = 64'h3636000000000000;
        font[8'h23] = 64'h36367F367F363600;
        font[8'h24] = 64'h0C3E031E301F0C00;
        font[8'h25] = 64'h006333180C666300;
        font[8'h26] = 64'h1C361C6E3B336E00;
        font[8'h27] = 64'h0606030000000000;
        font[8'h28] = 64'h180C0606060C1800;
        font[8'h29] = 64'h060C1818180C0600;
        font[8'h2a] = 64'h00663CFF3C660000;
        font[8'h2b] = 64'h000C0C3F0C0C0000;
        font[8'h2c] = 64'h00000000000C0C06;
        font[8'h2d] = 64'h0000003F00000000;
        font[8'h2e] = 64'h00000000000C0C00;
        font[8'h2f] = 64'h6030180C06030100;
        font[8'h30] = 64'h3E63737B6F673E00;
        font[8'h31] = 64'h0C0E0C0C0C0C3F00;
        font[8'h32] = 64'h1E33301C06333F00;
        font[8'h33] = 64'h1E33301C30331E00;
        font[8'h34] = 64'h383C36337F307800;
        font[8'h35] = 64'h3F031F3030331E00;
        font[8'h36] = 64'h1C06031F33331E00;
        font[8'h37] = 64'h3F3330180C0C0C00;
        font[8'h38] = 64'h1E33331E33331E00;
        font[8'h39] = 64'h1E33333E30180E00;
        font[8'h3a] = 64'h000C0C00000C0C00;
        font[8'h3b] = 64'h000C0C00000C0C06;
        font[8'h3c] = 64'h180C0603060C1800;
        font[8'h3d] = 64'h00003F00003F0000;
        font[8'h3e] = 64'h060C1830180C0600;
        font[8'h3f] = 64'h1E3330180C000C00;
        font[8'h40] = 64'h3E637B7B7B031E00;
        font[8'h41] = 64'h0C1E33333F333300;
        font[8'h42] = 64'h3F66663E66663F00;
        font[8'h43] = 64'h3C66030303663C00;
        font[8'h44] = 64'h1F36666666361F00;
        font[8'h45] = 64'h7F46161E16467F00;
        font[8'h46] = 64'h7F46161E16060F00;
        font[8'h47] = 64'h3C66030373667C00;
        font[8'h48] = 64'h3333333F33333300;
        font[8'h49] = 64'h1E0C0C0C0C0C1E00;
        font[8'h4a] = 64'h7830303033331E00;
        font[8'h4b] = 64'h6766361E36666700;
        font[8'h4c] = 64'h0F06060646667F00;
        font[8'h4d] = 64'h63777F7F6B636300;
        font[8'h4e] = 64'h63676F7B73636300;
        font[8'h4f] = 64'h1C36636363361C00;
        font[8'h50] = 64'h3F66663E06060F00;
        font[8'h51] = 64'h1E3333333B1E3800;
        font[8'h52] = 64'h3F66663E36666700;
        font[8'h53] = 64'h1E33070E38331E00;
        font[8'h54] = 64'h3F2D0C0C0C0C1E00;
        font[8'h55] = 64'h3333333333333F00;
        font[8'h56] = 64'h33333333331E0C00;
        font[8'h57] = 64'h6363636B7F776300;
        font[8'h58] = 64'h6363361C1C366300;
        font[8'h59] = 64'h3333331E0C0C1E00;
        font[8'h5a] = 64'h7F6331184C667F00;
        font[8'h5b] = 64'h1E06060606061E00;
        font[8'h5c] = 64'h03060C1830604000;
        font[8'h5d] = 64'h1E18181818181E00;
        font[8'h5e] = 64'h081C366300000000;
        font[8'h5f] = 64'h00000000000000FF;
        font[8'h60] = 64'h0C0C180000000000;
        font[8'h61] = 64'h00001E303E336E00;
        font[8'h62] = 64'h0706063E66663B00;
        font[8'h63] = 64'h00001E3303331E00;
        font[8'h64] = 64'h3830303e33336E00;
        font[8'h65] = 64'h00001E333f031E00;
        font[8'h66] = 64'h1C36060f06060F00;
        font[8'h67] = 64'h00006E33333E301F;
        font[8'h68] = 64'h0706366E66666700;
        font[8'h69] = 64'h0C000E0C0C0C1E00;
        font[8'h6a] = 64'h300030303033331E;
        font[8'h6b] = 64'h070666361E366700;
        font[8'h6c] = 64'h0E0C0C0C0C0C1E00;
        font[8'h6d] = 64'h0000337F7F6B6300;
        font[8'h6e] = 64'h00001F3333333300;
        font[8'h6f] = 64'h00001E3333331E00;
        font[8'h70] = 64'h00003B66663E060F;
        font[8'h71] = 64'h00006E33333E3078;
        font[8'h72] = 64'h00003B6E66060F00;
        font[8'h73] = 64'h00003E031E301F00;
        font[8'h74] = 64'h080C3E0C0C2C1800;
        font[8'h75] = 64'h0000333333336E00;
        font[8'h76] = 64'h00003333331E0C00;
        font[8'h77] = 64'h0000636B7F7F3600;
        font[8'h78] = 64'h000063361C366300;
        font[8'h79] = 64'h00003333333E301F;
        font[8'h7a] = 64'h00003F190C263F00;
        font[8'h7b] = 64'h380C0C070C0C3800;
        font[8'h7c] = 64'h1818180018181800;
        font[8'h7d] = 64'h070C0C380C0C0700;
        font[8'h7e] = 64'h6E3B000000000000;
        font[8'h7f] = 64'h0000000000000000;
    end

    always @ (posedge clk) bitmap <= ch[7] ? 64'h0000000000000000 : font[ch[6:0]];
endmodule
