module arp (
    input clk, input rst,
    output request, input grant,
    output valid, output error, output [7:0] data,
);
    
endmodule
